library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tt_um_top is
    port (
        ui_in1   : in  std_logic_vector(7 downto 0);
        ui_in2   : in  std_logic_vector(7 downto 0);
        ui_in3   : in  std_logic_vector(7 downto 0);
        
        uo_out1  : out std_logic_vector(7 downto 0);
        uo_out2  : out std_logic_vector(7 downto 0);
        uo_out3  : out std_logic_vector(7 downto 0);
        uo_out4  : out std_logic_vector(7 downto 0);


        ena     : in  std_logic;
        clk     : in  std_logic;
        rst_n   : in  std_logic
    );
end tt_um_top;


    
architecture Behavioral of tt_um_top is

 component boot_loader port (  rst : IN STD_LOGIC;
        clk : IN STD_LOGIC;
        ce : IN STD_LOGIC;
        rx : IN STD_LOGIC;
        tx : OUT STD_LOGIC;
        boot : OUT STD_LOGIC;
        scan_memory : IN STD_LOGIC;
        ram_out : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        ram_rw : OUT STD_LOGIC;
        ram_enable : OUT STD_LOGIC;
        ram_adr : OUT STD_LOGIC_VECTOR(RAM_ADR_WIDTH - 1 DOWNTO 0);
        ram_in : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
 end component ;

begin

   -- uo_out <= std_logic_vector(unsigned(ui_in) + unsigned(uio_in));
    uio_out <= "00000000";
    uio_oe <= "00000000";
    
     U1 : compteur  port map (
                            clk => clk,
                            rst => not(rst_n),
                            cmpt =>   uo_out
                        );


end Behavioral;
